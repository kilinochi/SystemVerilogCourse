`timescale 1 ns/ 100 ps
module b27s(sw, ss_a);
localparam N = 4;

(* altera_attribute = "-name IO_STANDARD \"3.3-V LVCMOS\"", chip_pin = "AF10, AF9, AC12, AB12" *)
input 			[N - 1:0]	sw;
(* altera_attribute = "-name IO_STANDARD \"3.3-V LVCMOS\"", chip_pin = "AH28, AG28, AF28, AG27, AE28, AE27, AE26" *)
output reg 		[2*N - 2:0]	ss_a;

reg			[6:0]		ss_arr	[15:0];

initial 
begin
	ss_arr[0]  = 7'h40; // 0
	ss_arr[1]  = 7'h79; // 1
	ss_arr[2]  = 7'h24; // 2
	ss_arr[3]  = 7'h30; // 3
	ss_arr[4]  = 7'h19; // 4
	ss_arr[5]  = 7'h12; // 5
	ss_arr[6]  = 7'h02; // 6
	ss_arr[7]  = 7'h78; // 7
	ss_arr[8]  = 7'h00; // 8
	ss_arr[9]  = 7'h10; // 9
	ss_arr[10] = 7'h08; // 10
	ss_arr[11] = 7'h03; // A
	ss_arr[12] = 7'h46; // B
	ss_arr[13] = 7'h21; // C
	ss_arr[14] = 7'h06; // D
	ss_arr[15] = 7'h0e; // F
end
	
always @*
begin
	ss_a = ss_arr[sw[N - 1:0]];
end

endmodule
